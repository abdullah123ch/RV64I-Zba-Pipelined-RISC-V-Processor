module decode (
    input  logic        clk,
    input  logic        rst,
    
    // Inputs from IF/ID Register
    input  logic [31:0] Instr_D,
    input  logic [63:0] PC_D,
    
    // Inputs from Writeback Stage (Feedback)
    input  logic [63:0] Result_W,    // Data to be written
    input  logic [4:0]  Rd_W,        // Destination register address
    input  logic        RegWrite_W,  // Write enable signal
    
    // Control Signals (To be generated by Controller)
    input  logic [2:0]  ImmSrc_D,    // For ImmGen
    
    // Outputs to ID/EX Register
    output logic [63:0] RD1_D,       // Register operand 1
    output logic [63:0] RD2_D,       // Register operand 2
    output logic [63:0] ImmExt_D,    // Sign-extended immediate
    output logic [4:0]  Rd_D,        // Destination register address
    output logic [63:0] PC_D_out     // Pass-through PC
);

    // 1. Internal wire for destination register extraction
    assign Rd_D = Instr_D[11:7];
    assign PC_D_out = PC_D;

    // 2. Instantiate Register File
    // Note: WD3 and A3 come from the Writeback (W) stage
    register rf (
        .clk(clk),
        .rst(rst),
        .A1(Instr_D[19:15]), // rs1
        .A2(Instr_D[24:20]), // rs2
        .A3(Rd_W),           // rd from WB stage
        .WD3(Result_W),      // data from WB stage
        .WE3(RegWrite_W),
        .RD1(RD1_D),
        .RD2(RD2_D)
    );

    // 3. Instantiate Immediate Generator
    immediate ig (
        .Instr(Instr_D),
        .ImmSrc(ImmSrc_D),
        .ImmExt(ImmExt_D)
    );

endmodule